module xx_regfile(

input   clk ,
input   rstn,
input   en  ,
input   we  ,
input   [31:0]  addr,
input   [31:0]  datai,
outupt wire  [31:0]  datao,
// regfile0

// regfile1

);
    
endmodule //xx_regfile
