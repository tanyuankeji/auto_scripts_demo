wire spi_clk_buf;
wire sclk_in;
wire spi_clk_n_0;
